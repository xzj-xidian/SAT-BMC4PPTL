/////////////////////////////////////////////////////////////////////
////                                                             ////
////  DES                                                        ////
////  DES Top Level module                                       ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2001 Rudolf Usselmann                         ////
////                    rudi@asics.ws                            ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////

module des(desOut, desIn, key, decrypt, roundSel, clk);
output	[63:0]	desOut;
input	[63:0]	desIn;
input	[55:0]	key;
input		decrypt;
input	[3:0]	roundSel;
input		clk;

wire	[1:48]	K_sub;
wire	[1:64]	IP, FP;
reg	[1:32]	L, R;
wire	[1:32]	Xin;
wire	[1:32]	Lout, Rout;
wire	[1:32]	out;

assign Lout = (roundSel == 0) ? IP[33:64] : R;
assign Xin  = (roundSel == 0) ? IP[01:32] : L;
assign Rout = Xin ^ out;
assign FP = { Rout, Lout};

crp u0( .P(out), .R(Lout), .K_sub(K_sub) );

always @(posedge clk)
        L <= #1 Lout;

always @(posedge clk)
        R <= #1 Rout;

// Select a subkey from key.
key_sel u1(
	.K_sub(		K_sub		),
	.K(		key		),
	.roundSel(	roundSel	),
	.decrypt(	decrypt		)
	);

// Perform initial permutation
assign IP[1:64] = {	desIn[06], desIn[14], desIn[22], desIn[30], desIn[38], desIn[46],
			desIn[54], desIn[62], desIn[04], desIn[12], desIn[20], desIn[28],
			desIn[36], desIn[44], desIn[52], desIn[60], desIn[02], desIn[10],
			desIn[18], desIn[26], desIn[34], desIn[42], desIn[50], desIn[58],
			desIn[00], desIn[08], desIn[16], desIn[24], desIn[32], desIn[40],
			desIn[48], desIn[56], desIn[07], desIn[15], desIn[23], desIn[31],
			desIn[39], desIn[47], desIn[55], desIn[63], desIn[05], desIn[13],
			desIn[21], desIn[29], desIn[37], desIn[45], desIn[53], desIn[61],
			desIn[03], desIn[11], desIn[19], desIn[27], desIn[35], desIn[43],
			desIn[51], desIn[59], desIn[01], desIn[09], desIn[17], desIn[25],
			desIn[33], desIn[41], desIn[49], desIn[57]};

// Perform final permutation
assign desOut = {	FP[40], FP[08], FP[48], FP[16], FP[56], FP[24], FP[64], FP[32],
			FP[39], FP[07], FP[47], FP[15], FP[55], FP[23], FP[63], FP[31],
			FP[38], FP[06], FP[46], FP[14], FP[54], FP[22], FP[62], FP[30],
			FP[37], FP[05], FP[45], FP[13], FP[53], FP[21], FP[61], FP[29],
			FP[36], FP[04], FP[44], FP[12], FP[52], FP[20], FP[60], FP[28],
			FP[35], FP[03], FP[43], FP[11], FP[51], FP[19], FP[59], FP[27],
			FP[34], FP[02], FP[42], FP[10], FP[50], FP[18], FP[58], FP[26],
			FP[33], FP[01], FP[41], FP[09], FP[49], FP[17], FP[57], FP[25] };

//p1: assert property (@(posedge clock) (roundSel != 0) |->  Lout == IP[33:64] && Xin = IP[01:32]);

//p2: assert property (@(posedge clock)  (R != 0) |-> (out != 0));

p3: assert property (@(posedge clock) ##[0:$] (desOut[0] == FP[40] && desOut[63] == FP[25]));

endmodule

module  crp(P, R, K_sub);
output	[1:32]	P;
input	[1:32]	R;
input	[1:48]	K_sub;

wire	[1:48] E;
wire	[1:48] X;
wire	[1:32] S;

assign E[1:48] = {	R[32], R[1], R[2], R[3], R[4], R[5], R[4], R[5],
			R[6], R[7], R[8], R[9], R[8], R[9], R[10], R[11],
			R[12], R[13], R[12], R[13], R[14], R[15], R[16],
			R[17], R[16], R[17], R[18], R[19], R[20], R[21],
			R[20], R[21], R[22], R[23], R[24], R[25], R[24],
			R[25], R[26], R[27], R[28], R[29], R[28], R[29],
			R[30], R[31], R[32], R[1]};

assign X = E ^ K_sub;

sbox1 u0( .addr(X[01:06]), .dout(S[01:04]) );
sbox2 u1( .addr(X[07:12]), .dout(S[05:08]) );
sbox3 u2( .addr(X[13:18]), .dout(S[09:12]) );
sbox4 u3( .addr(X[19:24]), .dout(S[13:16]) );
sbox5 u4( .addr(X[25:30]), .dout(S[17:20]) );
sbox6 u5( .addr(X[31:36]), .dout(S[21:24]) );
sbox7 u6( .addr(X[37:42]), .dout(S[25:28]) );
sbox8 u7( .addr(X[43:48]), .dout(S[29:32]) );

assign P[1:32] = {	S[16], S[7], S[20], S[21], S[29], S[12], S[28],
			S[17], S[1], S[15], S[23], S[26], S[5], S[18],
			S[31], S[10], S[2], S[8], S[24], S[14], S[32],
			S[27], S[3], S[9], S[19], S[13], S[30], S[6],
			S[22], S[11], S[4], S[25]};

endmodule


module  sbox1(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout =  14;
         1:  dout =   4;
         2:  dout =  13;
         3:  dout =   1;
         4:  dout =   2;
         5:  dout =  15;
         6:  dout =  11;
         7:  dout =   8;
         8:  dout =   3;
         9:  dout =  10;
        10:  dout =   6;
        11:  dout =  12;
        12:  dout =   5;
        13:  dout =   9;
        14:  dout =   0;
        15:  dout =   7;

        16:  dout =   0;
        17:  dout =  15;
        18:  dout =   7;
        19:  dout =   4;
        20:  dout =  14;
        21:  dout =   2;
        22:  dout =  13;
        23:  dout =   1;
        24:  dout =  10;
        25:  dout =   6;
        26:  dout =  12;
        27:  dout =  11;
        28:  dout =   9;
        29:  dout =   5;
        30:  dout =   3;
        31:  dout =   8;

        32:  dout =   4;
        33:  dout =   1;
        34:  dout =  14;
        35:  dout =   8;
        36:  dout =  13;
        37:  dout =   6;
        38:  dout =   2;
        39:  dout =  11;
        40:  dout =  15;
        41:  dout =  12;
        42:  dout =   9;
        43:  dout =   7;
        44:  dout =   3;
        45:  dout =  10;
        46:  dout =   5;
        47:  dout =   0;

        48:  dout =  15;
        49:  dout =  12;
        50:  dout =   8;
        51:  dout =   2;
        52:  dout =   4;
        53:  dout =   9;
        54:  dout =   1;
        55:  dout =   7;
        56:  dout =   5;
        57:  dout =  11;
        58:  dout =   3;
        59:  dout =  14;
        60:  dout =  10;
        61:  dout =   0;
        62:  dout =   6;
        63:  dout =  13;

    endcase
    end

endmodule

module  sbox2(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout = 15;
         1:  dout =  1;
         2:  dout =  8;
         3:  dout = 14;
         4:  dout =  6;
         5:  dout = 11;
         6:  dout =  3;
         7:  dout =  4;
         8:  dout =  9;
         9:  dout =  7;
        10:  dout =  2;
        11:  dout = 13;
        12:  dout = 12;
        13:  dout =  0;
        14:  dout =  5;
        15:  dout = 10;

        16:  dout =  3;
        17:  dout = 13;
        18:  dout =  4;
        19:  dout =  7;
        20:  dout = 15;
        21:  dout =  2;
        22:  dout =  8;
        23:  dout = 14;
        24:  dout = 12;
        25:  dout =  0;
        26:  dout =  1;
        27:  dout = 10;
        28:  dout =  6;
        29:  dout =  9;
        30:  dout = 11;
        31:  dout =  5;

        32:  dout =  0;
        33:  dout = 14;
        34:  dout =  7;
        35:  dout = 11;
        36:  dout = 10;
        37:  dout =  4;
        38:  dout = 13;
        39:  dout =  1;
        40:  dout =  5;
        41:  dout =  8;
        42:  dout = 12;
        43:  dout =  6;
        44:  dout =  9;
        45:  dout =  3;
        46:  dout =  2;
        47:  dout = 15;

        48:  dout = 13;
        49:  dout =  8;
        50:  dout = 10;
        51:  dout =  1;
        52:  dout =  3;
        53:  dout = 15;
        54:  dout =  4;
        55:  dout =  2;
        56:  dout = 11;
        57:  dout =  6;
        58:  dout =  7;
        59:  dout = 12;
        60:  dout =  0;
        61:  dout =  5;
        62:  dout = 14;
        63:  dout =  9;

    endcase
    end

endmodule


module  sbox3(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout = 10;
         1:  dout =  0;
         2:  dout =  9;
         3:  dout = 14;
         4:  dout =  6;
         5:  dout =  3;
         6:  dout = 15;
         7:  dout =  5;
         8:  dout =  1;
         9:  dout = 13;
        10:  dout = 12;
        11:  dout =  7;
        12:  dout = 11;
        13:  dout =  4;
        14:  dout =  2;
        15:  dout =  8;

        16:  dout = 13;
        17:  dout =  7;
        18:  dout =  0;
        19:  dout =  9;
        20:  dout =  3;
        21:  dout =  4;
        22:  dout =  6;
        23:  dout = 10;
        24:  dout =  2;
        25:  dout =  8;
        26:  dout =  5;
        27:  dout = 14;
        28:  dout = 12;
        29:  dout = 11;
        30:  dout = 15;
        31:  dout =  1;

        32:  dout = 13;
        33:  dout =  6;
        34:  dout =  4;
        35:  dout =  9;
        36:  dout =  8;
        37:  dout = 15;
        38:  dout =  3;
        39:  dout =  0;
        40:  dout = 11;
        41:  dout =  1;
        42:  dout =  2;
        43:  dout = 12;
        44:  dout =  5;
        45:  dout = 10;
        46:  dout = 14;
        47:  dout =  7;

        48:  dout =  1;
        49:  dout = 10;
        50:  dout = 13;
        51:  dout =  0;
        52:  dout =  6;
        53:  dout =  9;
        54:  dout =  8;
        55:  dout =  7;
        56:  dout =  4;
        57:  dout = 15;
        58:  dout = 14;
        59:  dout =  3;
        60:  dout = 11;
        61:  dout =  5;
        62:  dout =  2;
        63:  dout = 12;

    endcase
    end

endmodule


module  sbox4(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout =  7;
         1:  dout = 13;
         2:  dout = 14;
         3:  dout =  3;
         4:  dout =  0;
         5:  dout =  6;
         6:  dout =  9;
         7:  dout = 10;
         8:  dout =  1;
         9:  dout =  2;
        10:  dout =  8;
        11:  dout =  5;
        12:  dout = 11;
        13:  dout = 12;
        14:  dout =  4;
        15:  dout = 15;

        16:  dout = 13;
        17:  dout =  8;
        18:  dout = 11;
        19:  dout =  5;
        20:  dout =  6;
        21:  dout = 15;
        22:  dout =  0;
        23:  dout =  3;
        24:  dout =  4;
        25:  dout =  7;
        26:  dout =  2;
        27:  dout = 12;
        28:  dout =  1;
        29:  dout = 10;
        30:  dout = 14;
        31:  dout =  9;

        32:  dout = 10;
        33:  dout =  6;
        34:  dout =  9;
        35:  dout =  0;
        36:  dout = 12;
        37:  dout = 11;
        38:  dout =  7;
        39:  dout = 13;
        40:  dout = 15;
        41:  dout =  1;
        42:  dout =  3;
        43:  dout = 14;
        44:  dout =  5;
        45:  dout =  2;
        46:  dout =  8;
        47:  dout =  4;

        48:  dout =  3;
        49:  dout = 15;
        50:  dout =  0;
        51:  dout =  6;
        52:  dout = 10;
        53:  dout =  1;
        54:  dout = 13;
        55:  dout =  8;
        56:  dout =  9;
        57:  dout =  4;
        58:  dout =  5;
        59:  dout = 11;
        60:  dout = 12;
        61:  dout =  7;
        62:  dout =  2;
        63:  dout = 14;

    endcase
    end

endmodule


module  sbox5(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout =  2;
         1:  dout = 12;
         2:  dout =  4;
         3:  dout =  1;
         4:  dout =  7;
         5:  dout = 10;
         6:  dout = 11;
         7:  dout =  6;
         8:  dout =  8;
         9:  dout =  5;
        10:  dout =  3;
        11:  dout = 15;
        12:  dout = 13;
        13:  dout =  0;
        14:  dout = 14;
        15:  dout =  9;

        16:  dout = 14;
        17:  dout = 11;
        18:  dout =  2;
        19:  dout = 12;
        20:  dout =  4;
        21:  dout =  7;
        22:  dout = 13;
        23:  dout =  1;
        24:  dout =  5;
        25:  dout =  0;
        26:  dout = 15;
        27:  dout = 10;
        28:  dout =  3;
        29:  dout =  9;
        30:  dout =  8;
        31:  dout =  6;

        32:  dout =  4;
        33:  dout =  2;
        34:  dout =  1;
        35:  dout = 11;
        36:  dout = 10;
        37:  dout = 13;
        38:  dout =  7;
        39:  dout =  8;
        40:  dout = 15;
        41:  dout =  9;
        42:  dout = 12;
        43:  dout =  5;
        44:  dout =  6;
        45:  dout =  3;
        46:  dout =  0;
        47:  dout = 14;

        48:  dout = 11;
        49:  dout =  8;
        50:  dout = 12;
        51:  dout =  7;
        52:  dout =  1;
        53:  dout = 14;
        54:  dout =  2;
        55:  dout = 13;
        56:  dout =  6;
        57:  dout = 15;
        58:  dout =  0;
        59:  dout =  9;
        60:  dout = 10;
        61:  dout =  4;
        62:  dout =  5;
        63:  dout =  3;

    endcase
    end

endmodule


module  sbox6(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout = 12;
         1:  dout =  1;
         2:  dout = 10;
         3:  dout = 15;
         4:  dout =  9;
         5:  dout =  2;
         6:  dout =  6;
         7:  dout =  8;
         8:  dout =  0;
         9:  dout = 13;
        10:  dout =  3;
        11:  dout =  4;
        12:  dout = 14;
        13:  dout =  7;
        14:  dout =  5;
        15:  dout = 11;

        16:  dout = 10;
        17:  dout = 15;
        18:  dout =  4;
        19:  dout =  2;
        20:  dout =  7;
        21:  dout = 12;
        22:  dout =  9;
        23:  dout =  5;
        24:  dout =  6;
        25:  dout =  1;
        26:  dout = 13;
        27:  dout = 14;
        28:  dout =  0;
        29:  dout = 11;
        30:  dout =  3;
        31:  dout =  8;

        32:  dout =  9;
        33:  dout = 14;
        34:  dout = 15;
        35:  dout =  5;
        36:  dout =  2;
        37:  dout =  8;
        38:  dout = 12;
        39:  dout =  3;
        40:  dout =  7;
        41:  dout =  0;
        42:  dout =  4;
        43:  dout = 10;
        44:  dout =  1;
        45:  dout = 13;
        46:  dout = 11;
        47:  dout =  6;

        48:  dout =  4;
        49:  dout =  3;
        50:  dout =  2;
        51:  dout = 12;
        52:  dout =  9;
        53:  dout =  5;
        54:  dout = 15;
        55:  dout = 10;
        56:  dout = 11;
        57:  dout = 14;
        58:  dout =  1;
        59:  dout =  7;
        60:  dout =  6;
        61:  dout =  0;
        62:  dout =  8;
        63:  dout = 13;

    endcase
    end

endmodule


module  sbox7(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout =  4;
         1:  dout = 11;
         2:  dout =  2;
         3:  dout = 14;
         4:  dout = 15;
         5:  dout =  0;
         6:  dout =  8;
         7:  dout = 13;
         8:  dout =  3;
         9:  dout = 12;
        10:  dout =  9;
        11:  dout =  7;
        12:  dout =  5;
        13:  dout = 10;
        14:  dout =  6;
        15:  dout =  1;

        16:  dout = 13;
        17:  dout =  0;
        18:  dout = 11;
        19:  dout =  7;
        20:  dout =  4;
        21:  dout =  9;
        22:  dout =  1;
        23:  dout = 10;
        24:  dout = 14;
        25:  dout =  3;
        26:  dout =  5;
        27:  dout = 12;
        28:  dout =  2;
        29:  dout = 15;
        30:  dout =  8;
        31:  dout =  6;

        32:  dout =  1;
        33:  dout =  4;
        34:  dout = 11;
        35:  dout = 13;
        36:  dout = 12;
        37:  dout =  3;
        38:  dout =  7;
        39:  dout = 14;
        40:  dout = 10;
        41:  dout = 15;
        42:  dout =  6;
        43:  dout =  8;
        44:  dout =  0;
        45:  dout =  5;
        46:  dout =  9;
        47:  dout =  2;

        48:  dout =  6;
        49:  dout = 11;
        50:  dout = 13;
        51:  dout =  8;
        52:  dout =  1;
        53:  dout =  4;
        54:  dout = 10;
        55:  dout =  7;
        56:  dout =  9;
        57:  dout =  5;
        58:  dout =  0;
        59:  dout = 15;
        60:  dout = 14;
        61:  dout =  2;
        62:  dout =  3;
        63:  dout = 12;

    endcase
    end

endmodule


module  sbox8(addr, dout);
input	[1:6] addr;
output	[1:4] dout;
reg	[1:4] dout;

always @(addr) begin
    case ({addr[1], addr[6], addr[2:5]})	//synopsys full_case parallel_case
         0:  dout = 13;
         1:  dout =  2;
         2:  dout =  8;
         3:  dout =  4;
         4:  dout =  6;
         5:  dout = 15;
         6:  dout = 11;
         7:  dout =  1;
         8:  dout = 10;
         9:  dout =  9;
        10:  dout =  3;
        11:  dout = 14;
        12:  dout =  5;
        13:  dout =  0;
        14:  dout = 12;
        15:  dout =  7;

        16:  dout =  1;
        17:  dout = 15;
        18:  dout = 13;
        19:  dout =  8;
        20:  dout = 10;
        21:  dout =  3;
        22:  dout =  7;
        23:  dout =  4;
        24:  dout = 12;
        25:  dout =  5;
        26:  dout =  6;
        27:  dout = 11;
        28:  dout =  0;
        29:  dout = 14;
        30:  dout =  9;
        31:  dout =  2;

        32:  dout =  7;
        33:  dout = 11;
        34:  dout =  4;
        35:  dout =  1;
        36:  dout =  9;
        37:  dout = 12;
        38:  dout = 14;
        39:  dout =  2;
        40:  dout =  0;
        41:  dout =  6;
        42:  dout = 10;
        43:  dout = 13;
        44:  dout = 15;
        45:  dout =  3;
        46:  dout =  5;
        47:  dout =  8;

        48:  dout =  2;
        49:  dout =  1;
        50:  dout = 14;
        51:  dout =  7;
        52:  dout =  4;
        53:  dout = 10;
        54:  dout =  8;
        55:  dout = 13;
        56:  dout = 15;
        57:  dout = 12;
        58:  dout =  9;
        59:  dout =  0;
        60:  dout =  3;
        61:  dout =  5;
        62:  dout =  6;
        63:  dout = 11;

    endcase
    end

endmodule


module  key_sel(K_sub, K, roundSel, decrypt);
output [1:48] K_sub;
input [55:0] K;
input [3:0] roundSel;
input   decrypt;

reg  [1:48] K_sub;
wire [1:48] K1, K2, K3, K4, K5, K6, K7, K8;

////  Modified: for about Half slices decreased
wire [2:0] roundSelH;  // ADD Sakamoto
wire   decryptH;  // ADD Sakamoto

assign roundSelH[2:0] = roundSel[3] ? (~roundSel[2:0]) : roundSel[2:0];
assign decryptH  = decrypt ^ roundSel[3];

always @(K1 or K2 or K3 or K4 or K5 or K6 or K7 or K8 or roundSelH)
    case (roundSelH)    // synopsys full_case parallel_case
            0:  K_sub = K1;
            1:  K_sub = K2;
            2:  K_sub = K3;
            3:  K_sub = K4;
            4:  K_sub = K5;
            5:  K_sub = K6;
            6:  K_sub = K7;
            7:  K_sub = K8;
    endcase


assign K8[1]  = decryptH ? K[6]  : K[24];
assign K8[2]  = decryptH ? K[27] : K[20];
assign K8[3]  = decryptH ? K[10] : K[3] ;
assign K8[4]  = decryptH ? K[19] : K[12];
assign K8[5]  = decryptH ? K[54] : K[47];
assign K8[6]  = decryptH ? K[25] : K[18];
assign K8[7]  = decryptH ? K[11] : K[4] ;
assign K8[8]  = decryptH ? K[47] : K[40];
assign K8[9]  = decryptH ? K[13] : K[6] ;
assign K8[10] = decryptH ? K[32] : K[25];
assign K8[11] = decryptH ? K[55] : K[48];
assign K8[12] = decryptH ? K[3]  : K[53];
assign K8[13] = decryptH ? K[12] : K[5] ;
assign K8[14] = decryptH ? K[41] : K[34];
assign K8[15] = decryptH ? K[17] : K[10];
assign K8[16] = decryptH ? K[18] : K[11];
assign K8[17] = decryptH ? K[33] : K[26];
assign K8[18] = decryptH ? K[46] : K[39];
assign K8[19] = decryptH ? K[20] : K[13];
assign K8[20] = decryptH ? K[39] : K[32];
assign K8[21] = decryptH ? K[40] : K[33];
assign K8[22] = decryptH ? K[48] : K[41];
assign K8[23] = decryptH ? K[24] : K[17];
assign K8[24] = decryptH ? K[4]  : K[54];
assign K8[25] = decryptH ? K[52] : K[45];
assign K8[26] = decryptH ? K[15] : K[8] ;
assign K8[27] = decryptH ? K[9]  : K[2] ;
assign K8[28] = decryptH ? K[51] : K[44];
assign K8[29] = decryptH ? K[35] : K[28];
assign K8[30] = decryptH ? K[36] : K[29];
assign K8[31] = decryptH ? K[2]  : K[50];
assign K8[32] = decryptH ? K[45] : K[38];
assign K8[33] = decryptH ? K[8]  : K[1] ;
assign K8[34] = decryptH ? K[21] : K[14];
assign K8[35] = decryptH ? K[23] : K[16];
assign K8[36] = decryptH ? K[42] : K[35];
assign K8[37] = decryptH ? K[14] : K[7] ;
assign K8[38] = decryptH ? K[49] : K[42];
assign K8[39] = decryptH ? K[38] : K[31];
assign K8[40] = decryptH ? K[43] : K[36];
assign K8[41] = decryptH ? K[30] : K[23];
assign K8[42] = decryptH ? K[22] : K[15];
assign K8[43] = decryptH ? K[28] : K[21];
assign K8[44] = decryptH ? K[0]  : K[52];
assign K8[45] = decryptH ? K[1]  : K[49];
assign K8[46] = decryptH ? K[44] : K[37];
assign K8[47] = decryptH ? K[50] : K[43];
assign K8[48] = decryptH ? K[16] : K[9] ;

assign K7[1]  = decryptH ? K[20] : K[10];
assign K7[2]  = decryptH ? K[41] : K[6] ;
assign K7[3]  = decryptH ? K[24] : K[46];
assign K7[4]  = decryptH ? K[33] : K[55];
assign K7[5]  = decryptH ? K[11] : K[33];
assign K7[6]  = decryptH ? K[39] : K[4] ;
assign K7[7]  = decryptH ? K[25] : K[47];
assign K7[8]  = decryptH ? K[4]  : K[26];
assign K7[9]  = decryptH ? K[27] : K[17];
assign K7[10] = decryptH ? K[46] : K[11];
assign K7[11] = decryptH ? K[12] : K[34];
assign K7[12] = decryptH ? K[17] : K[39];
assign K7[13] = decryptH ? K[26] : K[48];
assign K7[14] = decryptH ? K[55] : K[20];
assign K7[15] = decryptH ? K[6]  : K[53];
assign K7[16] = decryptH ? K[32] : K[54];
assign K7[17] = decryptH ? K[47] : K[12];
assign K7[18] = decryptH ? K[3]  : K[25];
assign K7[19] = decryptH ? K[34] : K[24];
assign K7[20] = decryptH ? K[53] : K[18];
assign K7[21] = decryptH ? K[54] : K[19];
assign K7[22] = decryptH ? K[5]  : K[27];
assign K7[23] = decryptH ? K[13] : K[3] ;
assign K7[24] = decryptH ? K[18] : K[40];
assign K7[25] = decryptH ? K[7]  : K[31];
assign K7[26] = decryptH ? K[29] : K[49];
assign K7[27] = decryptH ? K[23] : K[43];
assign K7[28] = decryptH ? K[38] : K[30];
assign K7[29] = decryptH ? K[49] : K[14];
assign K7[30] = decryptH ? K[50] : K[15];
assign K7[31] = decryptH ? K[16] : K[36];
assign K7[32] = decryptH ? K[0]  : K[51];
assign K7[33] = decryptH ? K[22] : K[42];
assign K7[34] = decryptH ? K[35] : K[0] ;
assign K7[35] = decryptH ? K[37] : K[2] ;
assign K7[36] = decryptH ? K[1]  : K[21];
assign K7[37] = decryptH ? K[28] : K[52];
assign K7[38] = decryptH ? K[8]  : K[28];
assign K7[39] = decryptH ? K[52] : K[44];
assign K7[40] = decryptH ? K[2]  : K[22];
assign K7[41] = decryptH ? K[44] : K[9] ;
assign K7[42] = decryptH ? K[36] : K[1] ;
assign K7[43] = decryptH ? K[42] : K[7] ;
assign K7[44] = decryptH ? K[14] : K[38];
assign K7[45] = decryptH ? K[15] : K[35];
assign K7[46] = decryptH ? K[31] : K[23];
assign K7[47] = decryptH ? K[9]  : K[29];
assign K7[48] = decryptH ? K[30] : K[50];

assign K6[1]  = decryptH ? K[34] : K[53];
assign K6[2]  = decryptH ? K[55] : K[17];
assign K6[3]  = decryptH ? K[13] : K[32];
assign K6[4]  = decryptH ? K[47] : K[41];
assign K6[5]  = decryptH ? K[25] : K[19];
assign K6[6]  = decryptH ? K[53] : K[47];
assign K6[7]  = decryptH ? K[39] : K[33];
assign K6[8]  = decryptH ? K[18] : K[12];
assign K6[9]  = decryptH ? K[41] : K[3] ;
assign K6[10] = decryptH ? K[3]  : K[54];
assign K6[11] = decryptH ? K[26] : K[20];
assign K6[12] = decryptH ? K[6]  : K[25];
assign K6[13] = decryptH ? K[40] : K[34];
assign K6[14] = decryptH ? K[12] : K[6] ;
assign K6[15] = decryptH ? K[20] : K[39];
assign K6[16] = decryptH ? K[46] : K[40];
assign K6[17] = decryptH ? K[4]  : K[55];
assign K6[18] = decryptH ? K[17] : K[11];
assign K6[19] = decryptH ? K[48] : K[10];
assign K6[20] = decryptH ? K[10] : K[4] ;
assign K6[21] = decryptH ? K[11] : K[5] ;
assign K6[22] = decryptH ? K[19] : K[13];
assign K6[23] = decryptH ? K[27] : K[46];
assign K6[24] = decryptH ? K[32] : K[26];
assign K6[25] = decryptH ? K[21] : K[44];
assign K6[26] = decryptH ? K[43] : K[35];
assign K6[27] = decryptH ? K[37] : K[29];
assign K6[28] = decryptH ? K[52] : K[16];
assign K6[29] = decryptH ? K[8]  : K[0] ;
assign K6[30] = decryptH ? K[9]  : K[1] ;
assign K6[31] = decryptH ? K[30] : K[22];
assign K6[32] = decryptH ? K[14] : K[37];
assign K6[33] = decryptH ? K[36] : K[28];
assign K6[34] = decryptH ? K[49] : K[45];
assign K6[35] = decryptH ? K[51] : K[43];
assign K6[36] = decryptH ? K[15] : K[7] ;
assign K6[37] = decryptH ? K[42] : K[38];
assign K6[38] = decryptH ? K[22] : K[14];
assign K6[39] = decryptH ? K[7]  : K[30];
assign K6[40] = decryptH ? K[16] : K[8] ;
assign K6[41] = decryptH ? K[31] : K[50];
assign K6[42] = decryptH ? K[50] : K[42];
assign K6[43] = decryptH ? K[1]  : K[52];
assign K6[44] = decryptH ? K[28] : K[51];
assign K6[45] = decryptH ? K[29] : K[21];
assign K6[46] = decryptH ? K[45] : K[9] ;
assign K6[47] = decryptH ? K[23] : K[15];
assign K6[48] = decryptH ? K[44] : K[36];

assign K5[1]  = decryptH ? K[48] : K[39];
assign K5[2]  = decryptH ? K[12] : K[3] ;
assign K5[3]  = decryptH ? K[27] : K[18];
assign K5[4]  = decryptH ? K[4]  : K[27];
assign K5[5]  = decryptH ? K[39] : K[5] ;
assign K5[6]  = decryptH ? K[10] : K[33];
assign K5[7]  = decryptH ? K[53] : K[19];
assign K5[8]  = decryptH ? K[32] : K[55];
assign K5[9]  = decryptH ? K[55] : K[46];
assign K5[10] = decryptH ? K[17] : K[40];
assign K5[11] = decryptH ? K[40] : K[6] ;
assign K5[12] = decryptH ? K[20] : K[11];
assign K5[13] = decryptH ? K[54] : K[20];
assign K5[14] = decryptH ? K[26] : K[17];
assign K5[15] = decryptH ? K[34] : K[25];
assign K5[16] = decryptH ? K[3]  : K[26];
assign K5[17] = decryptH ? K[18] : K[41];
assign K5[18] = decryptH ? K[6]  : K[54];
assign K5[19] = decryptH ? K[5]  : K[53];
assign K5[20] = decryptH ? K[24] : K[47];
assign K5[21] = decryptH ? K[25] : K[48];
assign K5[22] = decryptH ? K[33] : K[24];
assign K5[23] = decryptH ? K[41] : K[32];
assign K5[24] = decryptH ? K[46] : K[12];
assign K5[25] = decryptH ? K[35] : K[30];
assign K5[26] = decryptH ? K[2]  : K[21];
assign K5[27] = decryptH ? K[51] : K[15];
assign K5[28] = decryptH ? K[7]  : K[2] ;
assign K5[29] = decryptH ? K[22] : K[45];
assign K5[30] = decryptH ? K[23] : K[42];
assign K5[31] = decryptH ? K[44] : K[8] ;
assign K5[32] = decryptH ? K[28] : K[23];
assign K5[33] = decryptH ? K[50] : K[14];
assign K5[34] = decryptH ? K[8]  : K[31];
assign K5[35] = decryptH ? K[38] : K[29];
assign K5[36] = decryptH ? K[29] : K[52];
assign K5[37] = decryptH ? K[1]  : K[51];
assign K5[38] = decryptH ? K[36] : K[0] ;
assign K5[39] = decryptH ? K[21] : K[16];
assign K5[40] = decryptH ? K[30] : K[49];
assign K5[41] = decryptH ? K[45] : K[36];
assign K5[42] = decryptH ? K[9]  : K[28];
assign K5[43] = decryptH ? K[15] : K[38];
assign K5[44] = decryptH ? K[42] : K[37];
assign K5[45] = decryptH ? K[43] : K[7] ;
assign K5[46] = decryptH ? K[0]  : K[50];
assign K5[47] = decryptH ? K[37] : K[1] ;
assign K5[48] = decryptH ? K[31] : K[22];

assign K4[1]  = decryptH ? K[5]  : K[25];
assign K4[2]  = decryptH ? K[26] : K[46];
assign K4[3]  = decryptH ? K[41] : K[4] ;
assign K4[4]  = decryptH ? K[18] : K[13];
assign K4[5]  = decryptH ? K[53] : K[48];
assign K4[6]  = decryptH ? K[24] : K[19];
assign K4[7]  = decryptH ? K[10] : K[5] ;
assign K4[8]  = decryptH ? K[46] : K[41];
assign K4[9]  = decryptH ? K[12] : K[32];
assign K4[10] = decryptH ? K[6]  : K[26];
assign K4[11] = decryptH ? K[54] : K[17];
assign K4[12] = decryptH ? K[34] : K[54];
assign K4[13] = decryptH ? K[11] : K[6] ;
assign K4[14] = decryptH ? K[40] : K[3] ;
assign K4[15] = decryptH ? K[48] : K[11];
assign K4[16] = decryptH ? K[17] : K[12];
assign K4[17] = decryptH ? K[32] : K[27];
assign K4[18] = decryptH ? K[20] : K[40];
assign K4[19] = decryptH ? K[19] : K[39];
assign K4[20] = decryptH ? K[13] : K[33];
assign K4[21] = decryptH ? K[39] : K[34];
assign K4[22] = decryptH ? K[47] : K[10];
assign K4[23] = decryptH ? K[55] : K[18];
assign K4[24] = decryptH ? K[3]  : K[55];
assign K4[25] = decryptH ? K[49] : K[16];
assign K4[26] = decryptH ? K[16] : K[7] ;
assign K4[27] = decryptH ? K[38] : K[1] ;
assign K4[28] = decryptH ? K[21] : K[43];
assign K4[29] = decryptH ? K[36] : K[31];
assign K4[30] = decryptH ? K[37] : K[28];
assign K4[31] = decryptH ? K[31] : K[49];
assign K4[32] = decryptH ? K[42] : K[9] ;
assign K4[33] = decryptH ? K[9]  : K[0] ;
assign K4[34] = decryptH ? K[22] : K[44];
assign K4[35] = decryptH ? K[52] : K[15];
assign K4[36] = decryptH ? K[43] : K[38];
assign K4[37] = decryptH ? K[15] : K[37];
assign K4[38] = decryptH ? K[50] : K[45];
assign K4[39] = decryptH ? K[35] : K[2] ;
assign K4[40] = decryptH ? K[44] : K[35];
assign K4[41] = decryptH ? K[0]  : K[22];
assign K4[42] = decryptH ? K[23] : K[14];
assign K4[43] = decryptH ? K[29] : K[51];
assign K4[44] = decryptH ? K[1]  : K[23];
assign K4[45] = decryptH ? K[2]  : K[52];
assign K4[46] = decryptH ? K[14] : K[36];
assign K4[47] = decryptH ? K[51] : K[42];
assign K4[48] = decryptH ? K[45] : K[8] ;

assign K3[1]  = decryptH ? K[19] : K[11];
assign K3[2]  = decryptH ? K[40] : K[32];
assign K3[3]  = decryptH ? K[55] : K[47];
assign K3[4]  = decryptH ? K[32] : K[24];
assign K3[5]  = decryptH ? K[10] : K[34];
assign K3[6]  = decryptH ? K[13] : K[5] ;
assign K3[7]  = decryptH ? K[24] : K[48];
assign K3[8]  = decryptH ? K[3]  : K[27];
assign K3[9]  = decryptH ? K[26] : K[18];
assign K3[10] = decryptH ? K[20] : K[12];
assign K3[11] = decryptH ? K[11] : K[3] ;
assign K3[12] = decryptH ? K[48] : K[40];
assign K3[13] = decryptH ? K[25] : K[17];
assign K3[14] = decryptH ? K[54] : K[46];
assign K3[15] = decryptH ? K[5]  : K[54];
assign K3[16] = decryptH ? K[6]  : K[55];
assign K3[17] = decryptH ? K[46] : K[13];
assign K3[18] = decryptH ? K[34] : K[26];
assign K3[19] = decryptH ? K[33] : K[25];
assign K3[20] = decryptH ? K[27] : K[19];
assign K3[21] = decryptH ? K[53] : K[20];
assign K3[22] = decryptH ? K[4]  : K[53];
assign K3[23] = decryptH ? K[12] : K[4] ;
assign K3[24] = decryptH ? K[17] : K[41];
assign K3[25] = decryptH ? K[8]  : K[2] ;
assign K3[26] = decryptH ? K[30] : K[52];
assign K3[27] = decryptH ? K[52] : K[42];
assign K3[28] = decryptH ? K[35] : K[29];
assign K3[29] = decryptH ? K[50] : K[44];
assign K3[30] = decryptH ? K[51] : K[14];
assign K3[31] = decryptH ? K[45] : K[35];
assign K3[32] = decryptH ? K[1]  : K[50];
assign K3[33] = decryptH ? K[23] : K[45];
assign K3[34] = decryptH ? K[36] : K[30];
assign K3[35] = decryptH ? K[7]  : K[1] ;
assign K3[36] = decryptH ? K[2]  : K[51];
assign K3[37] = decryptH ? K[29] : K[23];
assign K3[38] = decryptH ? K[9]  : K[31];
assign K3[39] = decryptH ? K[49] : K[43];
assign K3[40] = decryptH ? K[31] : K[21];
assign K3[41] = decryptH ? K[14] : K[8] ;
assign K3[42] = decryptH ? K[37] : K[0] ;
assign K3[43] = decryptH ? K[43] : K[37];
assign K3[44] = decryptH ? K[15] : K[9] ;
assign K3[45] = decryptH ? K[16] : K[38];
assign K3[46] = decryptH ? K[28] : K[22];
assign K3[47] = decryptH ? K[38] : K[28];
assign K3[48] = decryptH ? K[0]  : K[49];

assign K2[1]  = decryptH ? K[33] : K[54];
assign K2[2]  = decryptH ? K[54] : K[18];
assign K2[3]  = decryptH ? K[12] : K[33];
assign K2[4]  = decryptH ? K[46] : K[10];
assign K2[5]  = decryptH ? K[24] : K[20];
assign K2[6]  = decryptH ? K[27] : K[48];
assign K2[7]  = decryptH ? K[13] : K[34];
assign K2[8]  = decryptH ? K[17] : K[13];
assign K2[9]  = decryptH ? K[40] : K[4] ;
assign K2[10] = decryptH ? K[34] : K[55];
assign K2[11] = decryptH ? K[25] : K[46];
assign K2[12] = decryptH ? K[5]  : K[26];
assign K2[13] = decryptH ? K[39] : K[3] ;
assign K2[14] = decryptH ? K[11] : K[32];
assign K2[15] = decryptH ? K[19] : K[40];
assign K2[16] = decryptH ? K[20] : K[41];
assign K2[17] = decryptH ? K[3]  : K[24];
assign K2[18] = decryptH ? K[48] : K[12];
assign K2[19] = decryptH ? K[47] : K[11];
assign K2[20] = decryptH ? K[41] : K[5] ;
assign K2[21] = decryptH ? K[10] : K[6] ;
assign K2[22] = decryptH ? K[18] : K[39];
assign K2[23] = decryptH ? K[26] : K[47];
assign K2[24] = decryptH ? K[6]  : K[27];
assign K2[25] = decryptH ? K[22] : K[43];
assign K2[26] = decryptH ? K[44] : K[38];
assign K2[27] = decryptH ? K[7]  : K[28];
assign K2[28] = decryptH ? K[49] : K[15];
assign K2[29] = decryptH ? K[9]  : K[30];
assign K2[30] = decryptH ? K[38] : K[0] ;
assign K2[31] = decryptH ? K[0]  : K[21];
assign K2[32] = decryptH ? K[15] : K[36];
assign K2[33] = decryptH ? K[37] : K[31];
assign K2[34] = decryptH ? K[50] : K[16];
assign K2[35] = decryptH ? K[21] : K[42];
assign K2[36] = decryptH ? K[16] : K[37];
assign K2[37] = decryptH ? K[43] : K[9] ;
assign K2[38] = decryptH ? K[23] : K[44];
assign K2[39] = decryptH ? K[8]  : K[29];
assign K2[40] = decryptH ? K[45] : K[7] ;
assign K2[41] = decryptH ? K[28] : K[49];
assign K2[42] = decryptH ? K[51] : K[45];
assign K2[43] = decryptH ? K[2]  : K[23];
assign K2[44] = decryptH ? K[29] : K[50];
assign K2[45] = decryptH ? K[30] : K[51];
assign K2[46] = decryptH ? K[42] : K[8] ;
assign K2[47] = decryptH ? K[52] : K[14];
assign K2[48] = decryptH ? K[14] : K[35];

assign K1[1]  = decryptH ? K[40] : K[47];
assign K1[2]  = decryptH ? K[4]  : K[11];
assign K1[3]  = decryptH ? K[19] : K[26];
assign K1[4]  = decryptH ? K[53] : K[3] ;
assign K1[5]  = decryptH ? K[6]  : K[13];
assign K1[6]  = decryptH ? K[34] : K[41];
assign K1[7]  = decryptH ? K[20] : K[27];
assign K1[8]  = decryptH ? K[24] : K[6] ;
assign K1[9]  = decryptH ? K[47] : K[54];
assign K1[10] = decryptH ? K[41] : K[48];
assign K1[11] = decryptH ? K[32] : K[39];
assign K1[12] = decryptH ? K[12] : K[19];
assign K1[13] = decryptH ? K[46] : K[53];
assign K1[14] = decryptH ? K[18] : K[25];
assign K1[15] = decryptH ? K[26] : K[33];
assign K1[16] = decryptH ? K[27] : K[34];
assign K1[17] = decryptH ? K[10] : K[17];
assign K1[18] = decryptH ? K[55] : K[5] ;
assign K1[19] = decryptH ? K[54] : K[4] ;
assign K1[20] = decryptH ? K[48] : K[55];
assign K1[21] = decryptH ? K[17] : K[24];
assign K1[22] = decryptH ? K[25] : K[32];
assign K1[23] = decryptH ? K[33] : K[40];
assign K1[24] = decryptH ? K[13] : K[20];
assign K1[25] = decryptH ? K[29] : K[36];
assign K1[26] = decryptH ? K[51] : K[31];
assign K1[27] = decryptH ? K[14] : K[21];
assign K1[28] = decryptH ? K[1]  : K[8] ;
assign K1[29] = decryptH ? K[16] : K[23];
assign K1[30] = decryptH ? K[45] : K[52];
assign K1[31] = decryptH ? K[7]  : K[14];
assign K1[32] = decryptH ? K[22] : K[29];
assign K1[33] = decryptH ? K[44] : K[51];
assign K1[34] = decryptH ? K[2]  : K[9] ;
assign K1[35] = decryptH ? K[28] : K[35];
assign K1[36] = decryptH ? K[23] : K[30];
assign K1[37] = decryptH ? K[50] : K[2] ;
assign K1[38] = decryptH ? K[30] : K[37];
assign K1[39] = decryptH ? K[15] : K[22];
assign K1[40] = decryptH ? K[52] : K[0] ;
assign K1[41] = decryptH ? K[35] : K[42];
assign K1[42] = decryptH ? K[31] : K[38];
assign K1[43] = decryptH ? K[9]  : K[16];
assign K1[44] = decryptH ? K[36] : K[43];
assign K1[45] = decryptH ? K[37] : K[44];
assign K1[46] = decryptH ? K[49] : K[1] ;
assign K1[47] = decryptH ? K[0]  : K[7] ;
assign K1[48] = decryptH ? K[21] : K[28];

endmodule